/*
    cic_decimator_variable_ahb.v
    Variable Sample Rate CIC Decimator with AHB Interface

    Copyright 2021-2022 Hiryuu T. (PFMRLIB)

    Licensed under the Apache License, Version 2.0 (the "License");
    you may not use this file except in compliance with the License.
    You may obtain a copy of the License at

        http://www.apache.org/licenses/LICENSE-2.0

    Unless required by applicable law or agreed to in writing, software
    distributed under the License is distributed on an "AS IS" BASIS,
    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
    See the License for the specific language governing permissions and
    limitations under the License.
*/
module cic_decimator_varialble_ahb(
    // Clock and reset
    input  wire clk,
    input  wire reset_n,
    input  wire ce,

    // AXI-Stream I/O
    input  wire [15:0] tdata_s,
    input  wire        tvalid_s,
    output wire        tready_s,

    output reg  [15:0] tdata_m,
    output reg         tvalid_m,
    input  wire        tready_m,

    // AHB Control Interface
    // HCLK, HRESETn are combined into global signals.
    input  wire [31:0]     haddr_s,
    input  wire [2:0]      hburst_s,
    // Locked sequence (HMASTLOCK) is not used.
    // Protection option (HPROT[6:0]) is not used.
    input  wire [2:0]      hsize_s,
    // Secure transfer (HNONSEC) is not used.
    // Exclusive transfer (HEXCL) is not used.
    // Master identifier (HMASTER[3:0]) is not used.
    input  wire [1:0]      htrans_s,
    input  wire [31:0]     hwdata_s,
    input  wire            hwrite_s,

    output reg  [31:0]     hrdata_s,
    output reg  [31:0]     hreadyout_s,
    output reg             hresp_s,
    // Exlusive transfer is not available, thus HEXOKAY signal is not used.

    input  wire            hsel_s
);

	// Registers and fields
    // Control interface
    reg  [31:0] reg_ctrl;
    wire deci_enable = reg_ctrl[0];

    // LSB truncation of each stage
    reg  [31:0] reg_trunc_intg_0;
    reg  [31:0] reg_trunc_intg_1;

    wire [7:0] intg_trunc_0 = reg_trunc_intg_0[7:0];
    wire [7:0] intg_trunc_1 = reg_trunc_intg_0[15:8];
    wire [7:0] intg_trunc_2 = reg_trunc_intg_0[23:16];
    wire [7:0] intg_trunc_3 = reg_trunc_intg_0[31:24];
    wire [7:0] intg_trunc_4 = reg_trunc_intg_1[7:0];

    // Decimate ratio, only low 16 bit is available
    reg  [15:0] reg_dec_ratio;

    // Data input
	reg  [15:0] data_in;
	reg         data_valid;
	reg         proc_en;

	always @(posedge clk, negedge reset_n) begin
		if(!reset_n) begin
			data_in    <= 0;
			data_valid <= 1'b0;
			proc_en    <= 1'b0;
		end
		else begin
			if(tvalid_s && tready_s)
				data_in <= tdata_s;

			data_valid <= tvalid_s;
			proc_en    <= tready_m;
		end
	end

	assign tready_s = proc_en;

    // CIC_GENERATOR_BEGIN
    // Generated by Hogenaur Pruning Calculator
    // Time: 2022-9-30 11:48:29
    // Environment: Python 3.10.4 (tags/v3.10.4:9d38120, Mar 23 2022, 23:13:41) [MSC v.1929 64 bit (AMD64)] on win32
    wire signed [52:0] d_0;
    wire signed [46:0] d_1;
    wire signed [38:0] d_2;
    wire signed [31:0] d_3;
    wire signed [24:0] d_4;
    wire signed [23:0] d_5;
    wire signed [21:0] d_6;
    wire signed [20:0] d_7;
    wire signed [19:0] d_8;
    wire signed [19:0] d_9;

    integrator #(
    	.DW (53)
    ) intg_0(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && proc_en),

		.din  ({{37{tdata_s[15]}}, tdata_s}),
		.dout (d_0)
    );

    integrator #(
    	.DW (47)
    ) intg_1(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && proc_en),

		.din  (d_0 >>> intg_trunc_0),
		.dout (d_1)
    );

    integrator #(
    	.DW (39)
    ) intg_2(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && proc_en),

		.din  (d_1 >>> intg_trunc_1),
		.dout (d_2)
    );

    integrator #(
    	.DW (32)
    ) intg_3(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && proc_en),

		.din  (d_2 >>> intg_trunc_2),
		.dout (d_3)
    );

    integrator #(
    	.DW (25)
    ) intg_4(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && proc_en),

		.din  (d_3 >>> intg_trunc_3),
		.dout (d_4)
    );

    // Resample
    reg         [15:0] cycle;
    
    wire resample_en = (cycle == reg_dec_ratio - 1) && proc_en;

    always @(posedge clk, negedge reset_n) begin
        if(!reset_n)
            cycle <= 0;
        else begin
            if(cycle >= reg_dec_ratio - 1)
                cycle <= 0;
            else
                cycle <= cycle + 1;
        end
    end

    comb #(
    	.DW (24),
    	.M  (2)
    ) comb_0(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && resample_en),

		.din  (d_4 >>> intg_trunc_4),
		.dout (d_5)
    );

    comb #(
    	.DW (22),
    	.M  (2)
    ) comb_1(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && resample_en),

		.din  (d_5 >>> 1),
		.dout (d_6)
    );

    comb #(
    	.DW (21),
    	.M  (2)
    ) comb_2(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && resample_en),

		.din  (d_6 >>> 1),
		.dout (d_7)
    );

    comb #(
    	.DW (20),
    	.M  (2)
    ) comb_3(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && resample_en),

		.din  (d_7 >>> 1),
		.dout (d_8)
    );

    comb #(
    	.DW (20),
    	.M  (2)
    ) comb_4(
		.clk     (clk),
		.reset_n (reset_n),
		.ce      (ce && resample_en),

		.din  (d_8),
		.dout (d_9)
    );
  
    // CIC_GENERATOR_END

    // AXI-Stream output
	always @(*) begin
		if(deci_enable)
			tdata_m = d_9[19:4];
		else
			tdata_m = data_in;

		tvalid_m = resample_en;
	end

	`include "ahb_intf_cicdec.v"
endmodule