/*
    axis_sequencer.sv
    Sequencer of all AXI-Stream sequence

    Copyright 2021-2023 Hiryuu "Concordia" T. (PFMRLIB)

    Licensed under the Apache License, Version 2.0 (the "License");
    you may not use this file except in compliance with the License.
    You may obtain a copy of the License at

        http://www.apache.org/licenses/LICENSE-2.0

    Unless required by applicable law or agreed to in writing, software
    distributed under the License is distributed on an "AS IS" BASIS,
    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
    See the License for the specific language governing permissions and
    limitations under the License.
*/
`include "uvm_macros.svh"

class axis_sequencer extends uvm_sequencer;
    `uvm_component_utils(axis_sequencer)

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction
endclass